interface intf;
//input
logic signed [15:0] A, B;
logic [2:0] OP;//(operation code)
//output
logic signed [31:0] ALU_OUTPUT;

endinterface 
